//This document contains TestBench Code to Verify Single Core MESI L1 Cache specified in HAS3.0

hello there
